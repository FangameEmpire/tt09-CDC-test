module alu_Testbench();

endmodule // alu_Testbench
